<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>17.6394,19.25,82.8856,-13</PageViewport>
<gate>
<ID>2</ID>
<type>AA_MUX_2x1</type>
<position>41.5,12</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>16 </output>
<input>
<ID>SEL_0</ID>12 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>EE_VDD</type>
<position>37,9</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>8</ID>
<type>FF_GND</type>
<position>37,12</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>38,18</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>25.5,18</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>51.5,18</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>63.5,18</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_MUX_2x1</type>
<position>34,2.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>18 </output>
<input>
<ID>SEL_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>FF_GND</type>
<position>29.5,0.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_MUX_2x1</type>
<position>44.5,2.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>32 </output>
<input>
<ID>SEL_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>EE_VDD</type>
<position>40,4.5</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_MUX_2x1</type>
<position>54.5,6.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>23 </output>
<input>
<ID>SEL_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>34</ID>
<type>FF_GND</type>
<position>51,4.5</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_MUX_2x1</type>
<position>58.5,2</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>33 </output>
<input>
<ID>SEL_0</ID>23 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>EE_VDD</type>
<position>54.5,-0.5</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>40</ID>
<type>FF_GND</type>
<position>53.5,2</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_MUX_2x1</type>
<position>45,-5.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>28 </output>
<input>
<ID>SEL_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>EE_VDD</type>
<position>40,-5.5</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_MUX_2x1</type>
<position>64,-9.5</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>36 </output>
<input>
<ID>SEL_0</ID>28 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>EE_VDD</type>
<position>60,-12</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>52</ID>
<type>FF_GND</type>
<position>58.5,-10</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_MUX_2x1</type>
<position>64,-2</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>35 </output>
<input>
<ID>SEL_0</ID>32 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>FF_GND</type>
<position>59.5,-4</position>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_MUX_2x1</type>
<position>70.5,-6</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>37 </input>
<output>
<ID>OUT</ID>38 </output>
<input>
<ID>SEL_0</ID>35 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>60</ID>
<type>EE_VDD</type>
<position>67,-4</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>62</ID>
<type>GA_LED</type>
<position>75,-6</position>
<input>
<ID>N_in0</ID>38 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,13,39.5,13</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,10,37,11</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,11,39.5,11</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,14.5,41.5,18</points>
<connection>
<GID>2</GID>
<name>SEL_0</name></connection>
<intersection>15.5 2</intersection>
<intersection>18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,18,41.5,18</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41.5,15.5,54.5,15.5</points>
<intersection>41.5 0</intersection>
<intersection>54.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>54.5,9,54.5,15.5</points>
<connection>
<GID>32</GID>
<name>SEL_0</name></connection>
<intersection>15.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-3,28.5,18</points>
<intersection>-3 2</intersection>
<intersection>5 3</intersection>
<intersection>18 10</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-3,45,-3</points>
<connection>
<GID>42</GID>
<name>SEL_0</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>28.5,5,34,5</points>
<intersection>28.5 0</intersection>
<intersection>34 11</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>27.5,18,28.5,18</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>28.5 0</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>34,5,34,5</points>
<connection>
<GID>24</GID>
<name>SEL_0</name></connection>
<intersection>5 3</intersection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,4,38.5,11.5</points>
<intersection>4 1</intersection>
<intersection>11.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,4,38.5,4</points>
<intersection>32 8</intersection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38.5,11.5,43.5,11.5</points>
<intersection>38.5 0</intersection>
<intersection>43.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>43.5,11.5,43.5,12</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<intersection>11.5 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>32,3.5,32,4</points>
<intersection>3.5 9</intersection>
<intersection>4 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>32,3.5,32,3.5</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>32 8</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,1.5,32,1.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>29.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>29.5,1.5,29.5,1.5</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>1.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,5,44.5,5.5</points>
<connection>
<GID>28</GID>
<name>SEL_0</name></connection>
<intersection>5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,5.5,44.5,5.5</points>
<intersection>36 2</intersection>
<intersection>44.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>36,2.5,36,5.5</points>
<intersection>2.5 5</intersection>
<intersection>5.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>36,2.5,36,2.5</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>36 2</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,-0.5,48.5,16.5</points>
<intersection>-0.5 1</intersection>
<intersection>16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-0.5,48.5,-0.5</points>
<intersection>42.5 3</intersection>
<intersection>48.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,16.5,54.5,16.5</points>
<intersection>48.5 0</intersection>
<intersection>54.5 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>42.5,-6.5,42.5,1.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>-6.5 5</intersection>
<intersection>-0.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>42.5,-6.5,43,-6.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>42.5 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>54.5,16.5,54.5,18</points>
<intersection>16.5 2</intersection>
<intersection>18 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>53.5,18,54.5,18</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>54.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,3.5,42.5,3.5</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<connection>
<GID>28</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,11.5,59,16</points>
<intersection>11.5 1</intersection>
<intersection>16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,11.5,59,11.5</points>
<intersection>52.5 3</intersection>
<intersection>59 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59,16,65.5,16</points>
<intersection>59 0</intersection>
<intersection>65.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>52.5,7.5,52.5,11.5</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<intersection>11.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>65.5,16,65.5,18</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>16 2</intersection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51,5.5,52.5,5.5</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<connection>
<GID>32</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,4.5,58.5,6.5</points>
<connection>
<GID>36</GID>
<name>SEL_0</name></connection>
<intersection>6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,6.5,58.5,6.5</points>
<connection>
<GID>32</GID>
<name>OUT</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,0.5,54.5,1</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,1,56.5,1</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,3,56.5,3</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<connection>
<GID>36</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-4.5,43,-4.5</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<connection>
<GID>42</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47,-5.5,64,-5.5</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>64 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>64,-7,64,-5.5</points>
<connection>
<GID>46</GID>
<name>SEL_0</name></connection>
<intersection>-5.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-10.5,62,-10.5</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>60 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>60,-11,60,-10.5</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>-10.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-9,58.5,-8.5</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-8.5,62,-8.5</points>
<connection>
<GID>46</GID>
<name>IN_1</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,0.5,64,10</points>
<connection>
<GID>54</GID>
<name>SEL_0</name></connection>
<intersection>10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,10,64,10</points>
<intersection>46.5 2</intersection>
<intersection>64 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>46.5,2.5,46.5,10</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<intersection>10 1</intersection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-1,61,2</points>
<intersection>-1 1</intersection>
<intersection>2 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-1,62,-1</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>60.5,2,61,2</points>
<connection>
<GID>36</GID>
<name>OUT</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-3,62,-3</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<connection>
<GID>54</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-3.5,70.5,-2</points>
<connection>
<GID>58</GID>
<name>SEL_0</name></connection>
<intersection>-2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66,-2,70.5,-2</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<intersection>70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-9.5,67,-7</points>
<intersection>-9.5 2</intersection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67,-7,68.5,-7</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>67 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>66,-9.5,67,-9.5</points>
<connection>
<GID>46</GID>
<name>OUT</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>67,-5,68.5,-5</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<connection>
<GID>58</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72.5,-6,74,-6</points>
<connection>
<GID>62</GID>
<name>N_in0</name></connection>
<connection>
<GID>58</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>